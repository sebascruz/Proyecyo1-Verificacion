//////////////////////////////////////////////////////////////////////////////////////////////////////
//
// Deco.v
// 
// Este modulo sirve como Decodificador 
//
//////////////////////////////////////////////////////////////////////////////////////////////////////


module Deco (
    input WR,
    input [3:0] SEL, 
    output reg [11:0] WE
);
    
    always @(*) begin
        case ({WR, SEL})
            5'b10000 : WE = 12'b100000000000; //AL 
            5'b10001 : WE = 12'b010000000000; //CL
            5'b10010 : WE = 12'b001000000000; //DL
            5'b10011 : WE = 12'b000100000000; //BL
            5'b10100 : WE = 12'b000010000000; //AH
            5'b10101 : WE = 12'b000001000000; //CH
            5'b10110 : WE = 12'b100000100000; //DH
            5'b10111 : WE = 12'b100000010000; //BH
            5'b11000 : WE = 12'b100010000000; //AX
            5'b11001 : WE = 12'b010001000000; //CX
            5'b11010 : WE = 12'b001000100000; //DX
            5'b11011 : WE = 12'b000100010000; //BX
            5'b11100 : WE = 12'b000000001000; //SP
            5'b11101 : WE = 12'b000000000100; //BP
            5'b11110 : WE = 12'b000000000010; //SI
            5'b11111 : WE = 12'b000000000001; //DI

            default : WE = 12'b000000000000;  
        endcase
    end
endmodule