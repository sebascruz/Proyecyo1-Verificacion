//////////////////////////////////////////////////////////////////////////////////////////////////////
//
// Mux2x8.v
// 
// Este modulo sirve como Mux2x8
//
//////////////////////////////////////////////////////////////////////////////////////////////////////

module Mux2x8 (
    input [7:0] ENT1,
    input [7:0] ENT2,
    input SEL,
    output reg [7:0] OUT
);

always @(*) begin
    case (SEL)
        1'b0 : OUT = ENT1;
        1'b1 : OUT = ENT2; 
    endcase
end

endmodule